/* Automatically generated by meta-parse.py */

// Copyright (c) 2016, 2017 Massachusetts Institute of Technology

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

`include "ProcConfig.bsv"
`include "Opcodes.defines"

import RVTypes::*;

typedef struct {
    Maybe#(RegType) rs1;
    Maybe#(RegType) rs2;
    Maybe#(RegType) rs3;
    Maybe#(RegType) dst;
    ImmType imm;
} InstType deriving (Bits, Eq, FShow);

function InstType toInstType(Instruction inst);
    Maybe#(RegType) i = tagged Valid RtGpr;
    Maybe#(RegType) f = tagged Valid RtFpu;
    Maybe#(RegType) n = tagged Invalid;
    InstType ret = (case (inst) matches
            `LUI:           InstType{rs1: n, rs2: n, rs3: n, dst: i, imm: ItU   };
            `AUIPC:         InstType{rs1: n, rs2: n, rs3: n, dst: i, imm: ItU   };
            `JAL:           InstType{rs1: n, rs2: n, rs3: n, dst: i, imm: ItUJ  };
            `JALR:          InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `BEQ:           InstType{rs1: i, rs2: i, rs3: n, dst: n, imm: ItSB  };
            `BNE:           InstType{rs1: i, rs2: i, rs3: n, dst: n, imm: ItSB  };
            `BLT:           InstType{rs1: i, rs2: i, rs3: n, dst: n, imm: ItSB  };
            `BGE:           InstType{rs1: i, rs2: i, rs3: n, dst: n, imm: ItSB  };
            `BLTU:          InstType{rs1: i, rs2: i, rs3: n, dst: n, imm: ItSB  };
            `BGEU:          InstType{rs1: i, rs2: i, rs3: n, dst: n, imm: ItSB  };
            `LB:            InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `LH:            InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `LW:            InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `LBU:           InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `LHU:           InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `SB:            InstType{rs1: i, rs2: i, rs3: n, dst: n, imm: ItS   };
            `SH:            InstType{rs1: i, rs2: i, rs3: n, dst: n, imm: ItS   };
            `SW:            InstType{rs1: i, rs2: i, rs3: n, dst: n, imm: ItS   };
            `ADDI:          InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `SLTI:          InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `SLTIU:         InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `XORI:          InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `ORI:           InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `ANDI:          InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `ADD:           InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `SUB:           InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `SLL:           InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `SLT:           InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `SLTU:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `XOR:           InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `SRL:           InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `SRA:           InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `OR:            InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AND:           InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `FENCE:         InstType{rs1: n, rs2: n, rs3: n, dst: n, imm: ItNone};
            `FENCE_I:       InstType{rs1: n, rs2: n, rs3: n, dst: n, imm: ItNone};
            `LWU:           InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `LD:            InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `SD:            InstType{rs1: i, rs2: i, rs3: n, dst: n, imm: ItS   };
            `SLLI_32:       InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `SRLI_32:       InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `SRAI_32:       InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `SLLI_64:       InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `SRLI_64:       InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `SRAI_64:       InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `ADDIW:         InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `SLLIW:         InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `SRLIW:         InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `SRAIW:         InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItI   };
            `ADDW:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `SUBW:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `SLLW:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `SRLW:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `SRAW:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `MUL:           InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `MULH:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `MULHSU:        InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `MULHU:         InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `DIV:           InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `DIVU:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `REM:           InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `REMU:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `MULW:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `DIVW:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `DIVUW:         InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `REMW:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `REMUW:         InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `LR_W:          InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItNone};
            `SC_W:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOSWAP_W:     InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOADD_W:      InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOXOR_W:      InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOOR_W:       InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOAND_W:      InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOMIN_W:      InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOMAX_W:      InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOMINU_W:     InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOMAXU_W:     InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `LR_D:          InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItNone};
            `SC_D:          InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOSWAP_D:     InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOADD_D:      InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOXOR_D:      InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOOR_D:       InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOAND_D:      InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOMIN_D:      InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOMAX_D:      InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOMINU_D:     InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `AMOMAXU_D:     InstType{rs1: i, rs2: i, rs3: n, dst: i, imm: ItNone};
            `ECALL:         InstType{rs1: n, rs2: n, rs3: n, dst: n, imm: ItNone};
            `EBREAK:        InstType{rs1: n, rs2: n, rs3: n, dst: n, imm: ItNone};
            `URET:          InstType{rs1: n, rs2: n, rs3: n, dst: n, imm: ItNone};
            `SRET:          InstType{rs1: n, rs2: n, rs3: n, dst: n, imm: ItNone};
            `HRET:          InstType{rs1: n, rs2: n, rs3: n, dst: n, imm: ItNone};
            `MRET:          InstType{rs1: n, rs2: n, rs3: n, dst: n, imm: ItNone};
            `DRET:          InstType{rs1: n, rs2: n, rs3: n, dst: n, imm: ItNone};
            `SFENCE_VM:     InstType{rs1: i, rs2: n, rs3: n, dst: n, imm: ItNone};
            `WFI:           InstType{rs1: n, rs2: n, rs3: n, dst: n, imm: ItNone};
            `CSRRW:         InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItNone};
            `CSRRS:         InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItNone};
            `CSRRC:         InstType{rs1: i, rs2: n, rs3: n, dst: i, imm: ItNone};
            `CSRRWI:        InstType{rs1: n, rs2: n, rs3: n, dst: i, imm: ItZ   };
            `CSRRSI:        InstType{rs1: n, rs2: n, rs3: n, dst: i, imm: ItZ   };
            `CSRRCI:        InstType{rs1: n, rs2: n, rs3: n, dst: i, imm: ItZ   };
            `FLW:           InstType{rs1: i, rs2: n, rs3: n, dst: f, imm: ItI   };
            `FSW:           InstType{rs1: i, rs2: f, rs3: n, dst: n, imm: ItS   };
            `FMADD_S:       InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: ItNone};
            `FMSUB_S:       InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: ItNone};
            `FNMSUB_S:      InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: ItNone};
            `FNMADD_S:      InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: ItNone};
            `FADD_S:        InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FSUB_S:        InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FMUL_S:        InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FDIV_S:        InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FSGNJ_S:       InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FSGNJN_S:      InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FSGNJX_S:      InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FMIN_S:        InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FMAX_S:        InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FSQRT_S:       InstType{rs1: f, rs2: n, rs3: n, dst: f, imm: ItNone};
            `FLE_S:         InstType{rs1: f, rs2: f, rs3: n, dst: i, imm: ItNone};
            `FLT_S:         InstType{rs1: f, rs2: f, rs3: n, dst: i, imm: ItNone};
            `FEQ_S:         InstType{rs1: f, rs2: f, rs3: n, dst: i, imm: ItNone};
            `FCVT_W_S:      InstType{rs1: f, rs2: n, rs3: n, dst: i, imm: ItNone};
            `FCVT_WU_S:     InstType{rs1: f, rs2: n, rs3: n, dst: i, imm: ItNone};
            `FCVT_S_W:      InstType{rs1: i, rs2: n, rs3: n, dst: f, imm: ItNone};
            `FCVT_S_WU:     InstType{rs1: i, rs2: n, rs3: n, dst: f, imm: ItNone};
            `FMV_X_S:       InstType{rs1: f, rs2: n, rs3: n, dst: i, imm: ItNone};
            `FCLASS_S:      InstType{rs1: f, rs2: n, rs3: n, dst: i, imm: ItNone};
            `FMV_S_X:       InstType{rs1: i, rs2: n, rs3: n, dst: f, imm: ItNone};
            `FCVT_L_S:      InstType{rs1: f, rs2: n, rs3: n, dst: i, imm: ItNone};
            `FCVT_LU_S:     InstType{rs1: f, rs2: n, rs3: n, dst: i, imm: ItNone};
            `FCVT_S_L:      InstType{rs1: i, rs2: n, rs3: n, dst: f, imm: ItNone};
            `FCVT_S_LU:     InstType{rs1: i, rs2: n, rs3: n, dst: f, imm: ItNone};
            `FLD:           InstType{rs1: i, rs2: n, rs3: n, dst: f, imm: ItI   };
            `FSD:           InstType{rs1: i, rs2: f, rs3: n, dst: n, imm: ItS   };
            `FMADD_D:       InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: ItNone};
            `FMSUB_D:       InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: ItNone};
            `FNMSUB_D:      InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: ItNone};
            `FNMADD_D:      InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: ItNone};
            `FADD_D:        InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FSUB_D:        InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FMUL_D:        InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FDIV_D:        InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FSGNJ_D:       InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FSGNJN_D:      InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FSGNJX_D:      InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FMIN_D:        InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FMAX_D:        InstType{rs1: f, rs2: f, rs3: n, dst: f, imm: ItNone};
            `FCVT_S_D:      InstType{rs1: f, rs2: n, rs3: n, dst: f, imm: ItNone};
            `FCVT_D_S:      InstType{rs1: f, rs2: n, rs3: n, dst: f, imm: ItNone};
            `FSQRT_D:       InstType{rs1: f, rs2: n, rs3: n, dst: f, imm: ItNone};
            `FLE_D:         InstType{rs1: f, rs2: f, rs3: n, dst: i, imm: ItNone};
            `FLT_D:         InstType{rs1: f, rs2: f, rs3: n, dst: i, imm: ItNone};
            `FEQ_D:         InstType{rs1: f, rs2: f, rs3: n, dst: i, imm: ItNone};
            `FCVT_W_D:      InstType{rs1: f, rs2: n, rs3: n, dst: i, imm: ItNone};
            `FCVT_WU_D:     InstType{rs1: f, rs2: n, rs3: n, dst: i, imm: ItNone};
            `FCVT_D_W:      InstType{rs1: i, rs2: n, rs3: n, dst: f, imm: ItNone};
            `FCVT_D_WU:     InstType{rs1: i, rs2: n, rs3: n, dst: f, imm: ItNone};
            `FCLASS_D:      InstType{rs1: f, rs2: n, rs3: n, dst: i, imm: ItNone};
            `FCVT_L_D:      InstType{rs1: f, rs2: n, rs3: n, dst: i, imm: ItNone};
            `FCVT_LU_D:     InstType{rs1: f, rs2: n, rs3: n, dst: i, imm: ItNone};
            `FMV_X_D:       InstType{rs1: f, rs2: n, rs3: n, dst: i, imm: ItNone};
            `FCVT_D_L:      InstType{rs1: i, rs2: n, rs3: n, dst: f, imm: ItNone};
            `FCVT_D_LU:     InstType{rs1: i, rs2: n, rs3: n, dst: f, imm: ItNone};
            `FMV_D_X:       InstType{rs1: i, rs2: n, rs3: n, dst: f, imm: ItNone};
            default:        ?;
        endcase);
    if ((ret.dst == tagged Valid RtGpr) && (getInstFields(inst).rd == 0)) begin
        ret.dst = tagged Invalid;
    end
    return ret;
endfunction
